module BCD_to_xs3(b,x);
input [3:0]b;
output [3:0]x;
wire w,y;
not(x[0],b[0]);

xnor(x[1],b[1],b[0]);

or(w,b[1],b[0]);
xor(x[2],b[2],w);

and(y,b[2],w);
or(x[3],b[3],y);
endmodule

module TB_BX();
reg [3:0]b;
wire [3:0]x;
BCD_to_xs3 BX1(b,x);
initial begin
#0 b=4'd0;
#100 b=4'd1;
#100 b=4'd2;
#100 b=4'd3;
#100 b=4'd4;
#100 b=4'd5;
#100 b=4'd6;
#100 b=4'd7;
#100 b=4'd8;
#100 b=4'd9;
#100 b=4'd10;
#100 b=4'd11;
#100 b=4'd12;
#100 b=4'd13;
#100 b=4'd14;
#100 b=4'd15;
end
endmodule

